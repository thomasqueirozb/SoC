
module niosLab2 (
	clk_clk,
	reset_reset_n,
	leds_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[5:0]	leds_export;
endmodule
